library verilog;
use verilog.vl_types.all;
entity checkpoint2 is
end checkpoint2;
