library verilog;
use verilog.vl_types.all;
entity checkpoint1 is
end checkpoint1;
